module QR;initial begin $write("%s",("Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[write,format=\"\"%s%s%s%s\"\",\"& VbLf &\"(\"\"\\\\write{-}{txt}{(\\\"\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put_Line(\\\\\\\\\\\"\"print\\\\\\\\\\\"\"\\\\\\\\\\\"\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"2\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR160,c:=b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"8\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR165,t:=\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"write('implement main()=print(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"BEGIN\\\\{s=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"d=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"(a#include<stdio.h>!nint main()\\\\{puts(!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"&3dlaiostream>!!n(3f5astd::cout<<(!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"class Program\\\\{public static void M93a@aSystem.Console.Write(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"let f(c :Int):Latin1=if c=127then!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3craelse(string_of c@x3cma g caffeine s3cba@,3oea!!!!!!!!Z3dra)@f(c+1)in print(x3ctaQuine Relay Coffee.<3dmanIngredientsu3eja!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@f 10r4igaMethod*3i%a);let g(String ->[])!!!!!!!!n[c;t]->74idaPut05wpa(int_of_char c)k6euainto the mixing bowl44klag t!!!!!!!!n|_ #4ktaLiquify contents ofQ3qeaPour)3w54elabaking dishL6fiaServes 1H4jeain g94dea)))sk3b[2cca!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" [2bw3kparts(nltnirp(])]~3kja.NUR POTSx3k,3l!$3zba!!&4l!$3lJ4nda[))r3kq3mL3k!$3|[2\\\\{ca\\\\};F3Aka)1(f\\\\{#qp]\\\\}Q3Dfa3(f\\\\{#K3Bga7(f\\\\{#.L3Bca51>4Fba105Gga36(f\\\\{#\\\\}6Bra21(f\\\\{# D ; EYB RCb;|X3(da,43O3HdaDNEE4[O39da. A36[O3<eaPOTSF4[46=36[O3:maRQ margorp d6HeP4[O31baS;6[O3;A4[JC2ca52A4[A4<ba&m8[C49gaS POOLoA[O3<ea\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&,)F4[oA;ga. TNUO76[O3:fa(rahcr:[96<gaB OD 0rA[O3;ca&,C4[H=8ca)A|8[3?<eaTXENz8[z8=66[dJ=haROF PUDK4[jJ[A4[j:rwa;TIUQ;)s(maertSesolC;)#ZBX4Kla115(f\\\\{#n\\\\})2i3aL4[O32ca3608Ema3(f\\\\{#(tnirP;85Bda369+6[O37ia402(f\\\\{#\\\\}D4[a<3ka904(f\\\\{#mif!$7CK;Lda918L;cj3bM4[M42ca34N;[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'A;oa99(f\\\\"));
$write("%s",("{#;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\})426y:aS4[R35ea0603F4[?69da134XVaja,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(rt.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'m<[??5ba6@HF:6Nha933(f\\\\{#nL[:53ca83.6ahaq\\\\})2173:6[v::ca76H=F:6T!$8[oC4ca21t8[pC;1Oaca\\\\}\\\\}5H[x8[D4[%?pca17pJFw8Nea7667\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'?bba4:6c96[UM3VT[-Q<gLai:[N;;ea&dne==[.X5ba8@M[R3:ca25<5az8[gJ>da825LD[\\\\{A:ca58\\\\}Qa:6[)?3ba5/6[*?<ba7j:[)?@\\\\}a&&PUEVIGESAELPn&&&&1,TUODAERs3ak5[XM3ba8Q3a:8[XM6ba5NV[F?Cea6940;6[c>;ca85F?[5Q[D4[i:rca105Q[s8:da738F?b~a(etirw;\\\\};u=:c;))652%%)u-c((||M6[78[D4[MHnca72e<FnWOda011C?coW[,:;da592:6[Y=9da343k:[EJCda#-<I4[)U3ba4y8[UX:ba9IQay8[)?4ba4xUG*?Pba9)?[)?Dba13Q[*?<R;ak:[)?>da||ilJ[p:5ca69\\\\{8[B=:ca76\\\\{8[OVBea2727:6[%S:ba1%8FvQ[D4[|Z-ba7|H[s8:ca95vQala&&&#BUS1,OD96[#8[D4[?Moba2ZR[@M;ba1VKapJNh;[t9;h:[h:[h"));
$write("%s",("Z+\\\\}Xa!$7[iZ7ba2,?bta(etirw;)3/4%%i(&&&&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'RC8?[D4[O3+ca82rCa/8[MM5da905IV[N4Bda59896[:5:ca47j:[HVBgaESAELPL4[IV3ca46|8[IV:ca99|8[IVDba0,I[IV;ba3H5a:6[LD[D4[JVoba5KD[JV;ba7*Qa\\\\}JeQa\\\\}2=:/t;2%%t+2*u=:u\\\\{od7 ot0 yreve;i-=:u;1=:+i\\\\{od))1(evom(dro=:t elihw?s;)s*||-7[O32ca69B5a.7[#@5TUbY:[#@?ca368>Gk;Oda573#@[#@[D4[AWsca10t8[AW;ca26#@bha#-<1,OD86[~8[D4[BEpba7\\\\}8[BE;ba83W[F5Bda62596[R39da211j:[4WCgKbxZDN4Iea5962#8[D=:ca63#8[sJCca06*HF:6Nda720.?[C=9ba4~Q[vA<ba9j:[.?Cmbn&&&&dohtem dne.n&&&&nrutern&&&&V);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovnin&&&&R5[O34lDa\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'9[FW5ba5>Ga\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'9[FW?\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'Kb:6[UE6TNG&R[D4[<G,da136s8[s89ca700Yaba&[2aeb\\\\}\\\\}\\\\}\\\\};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]+"));
$write("%s",("+n[c;y:]q[c?n<q=y\\\\{)0>2%%++i(fi;48%%)31-)i:3c+as(+87*q=q\\\\{);)(htgnel.s<i;(rof;n)rahc(+l8[Q9[D4[Z@nba7zP[:5;ca07zPazY[1=>ba5yP[0=:ba3yPbj:[#84zP[Q;=zPaaAb[2c=6[2?[D4[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'8oba8zO[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'8<ca542?[N4Cca4996[%8:ca96j:[\\\\}YB[2goa=]n[c);621<n++;Jaqa0=q,0=n,0=i tni;\\\\{5[~E2ca95PO[iU;ca79J8[DXBea6524:6[%89ca31H5a:6[\\\\{E[D4[ZVoba7zE[0Z;ba6.LaV?jMc6a2b9a*I2a4a5azbud;axb+b.b2b/cvbGa6a2b5a:fLa4a/c@cQtyb4aJaJa:f-a?Xxbrfzc6a/a6aHb<b<bHa6a6a>a9a@a3a?a7a|bKaKao5:a@aEa2aCtub8aucSjrS/apdxfMt5amdfb@rfdbdZcXcVc1bTcpcQc>a>aBh|zwbP4+bwbRZ9b5-RZ8bLaJaKa8bSJ>a:aJaJa8bTa.ZJaJa:b:aLaJaHaJaJaLaJa8bpBNaP4\\\\}bu3a+a8bpBm=4b|z;a8bm=wbRZ5-RZ|z9bLaMa\\\\}bJaNaI3oea|zvf84agaP4+bvfU3eea|zwbm3c1aJa0HVa;aW7Ua:aUa:ad|/apd8bMb1btb-aXcvb-a1bTc46acawb[5a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'aBh"));
$write("%s",("1e6aTs>a3a6a\\\\}bft5aKaKaCtucSj*b*b46cma8aubJawupbCa66aCa\\\\}bUcScucSj/a-s6aEa9aucDh/a-sub8aub5a/bxb1bJawbpcQcHa6a/a-s3b5aH4imaUcSc6aub8aQc|4aK7a4a<bRcef1dHa:f;a/aIduc=u8aQc/aIdHb|c8azc6azb9a2b9w3beaSdQck3cka/apdxbvbm484acaHa13gbaS/3ddaSdS/3n=apboc+bwdudTanbJazbHa6a-e9a-e7a|b9a6aQc<b=a-a\\\\{tVcNe1b6a6ao3ada|b9i3fEard7apbPH,d*d|dzdnd?B3bofBe+bLrcc7aPH5a2b@rMa\\\\{tVcjevbJa>a2a:boc:hu3akaxbDbyb4c6a33kSaxb1btbPZ4c/aId=a=aIdRdlbOa-aRalbOakb7vXa5rGdEdggCrfe?a/f4r4a0ejf?lKfAr|b4b0b=s\\\\}3eeaMgJe-5aware>i-b<iceBuKrjbGale:cf>cbbPa;aBeld8bfbpbfeubFcWbvbB2nbfeyeicYeyejeo2/f4rEmEa?aMs=l7h\\\\}p>a9a7b2cye:z,b-b\\\\}p=a9a7bubxbs3e53gbaA53lG3a53gja,p:r9a7b+)3flaAaddBaTs7bw-3bmaa|XbP\\\\{;i-b\\\\}pi3auayexdvdtd-b3p5f-bko,rl6awa9dug6i0r\\\\}rzr;hgmzr-r.r*6ecaxp\\\\{3axa\\\\{rxr,rJe0e=ast;h1"));
$write("%s",("b4bNe1V6hca:q/3aca-rg3kU3gcakh\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'3qg3\\\\{G3amaJele:bKfAr9aS3acaHmS35g39faDh2a2*4bca\\\\}nt4[g3i+7ama>lkg:fDrafof%7aCa@a>a8a6afepb-fCrKf;hJarcJa7b4eReZcfe>lkgybdh>l:rJa6afe7b5aKfArM3aba0?3fwa9a9b9a@aCa>lkgYsCrfe>au3cba@u3fwa@a>a:a|b9a0b9a@a>a7a6aw3aoaIa|b4e:a9bJa0b73ch4a&a@aCa9aCaAaJa9b>lkgnbff|c6areSj>l:@:b@4e|a4eNttbye>anbfe9apbfe?akuioyQ9b17/DK[R39u9Aga*b.bbbp67,4Adaye7*4[S5!$*4[*4wqanbKfTjTeSQxb1b6a9;a=a8b9a7b4eMaJayb>a-+le>aJaVcvgquTc0e<breIeff|c,bD\\\\{>aJa-b-a\\\\}3ccaBre=c+a<a2b4e+b|bxbvb:a>a>arc4e+b*eo2,b4b-b\\\\{c\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'Cgca;mO5[g3oRHocayl|4[g3[g3\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'ka2raf-b\\\\}ejop4[g3[1;)!$8aca|iv4[g3[g3[g3[z8U6a;awbof6afeYPc1:Zxd5bxb;uessteu>uVrYr;u|ursDuiuBu2w3b>cCs,6gAzb/0CzBaUvDauD4YxVRa*dzbPWCz*dTvRvPvNvB80v5-TatUEaYvybOaK-l@,bB"));
$write("%s",("+4@RUBat*Aa4wEV<5R*rU.zr|cvD\\\\},?ivk*Xu,71b8PzxWac1:Z=aSaVaJUe|aC*bf,1U48*b3UybdbCvQP:W\\\\}B<5jbhb,b@W?V@v8A-9JUZw29pO7=Y+z,\\\\{FCYdNx8*dybzbV|kbm=\\\\}w<a?aYajbvbkbeL*bpSdb=s3bVba/vD@+Z4*y?/2b*T@+e>kTP,CaPH/ZP,Cv9blb3Ul.;5iz,bZ4a/e\\\\{8\\\\{mTgxUv|8z8j\\\\}fTdTPLxP6zjS=EcvSSSaa|Vujb>;4v3S2bUa\\\\{SBSSauT6;Yv?|uTkbm=7SmxdNxbhb48*bUaa,8vUZ|Scv==ST=\\\\{XX\\\\{OjbZacxi3e5a9a=Ei3,v,\\\\{CvAv0v7b6SAvevdbAaTRi3QRdbOvYaCa3b@aVAhbTAFW57abbfzoSE6lb0v*RZu6EzRS|c6-:*Yhb>|jRjDdyeRcRo5ZQqv:wD\\\\}hbQd|vTQJFJwJFZaOQqvtdIN\\\\{vjbOaNufQ=ajbw3aWa+b<aXLqv?QxE=?D;Wu=a3UhbVTB4Byo5T\\\\{K*hb,RByFwnD5wixDaed?QxEKIfxGvedr,pQg5mQdwv-3Kd|h4aOa=\\\\{XXmGbbcQFz?a;xu\\\\{8zlbKzBPHOqw3-F8lOYH3Sk+e\\\\}VxaUYOmYZObw-DQxi\\\\{12E6gxiP30uv33gAaqwlbF?v,7=UUPLPBabd/,b?\\\\{F8wxBVaD4.JzfYBV\\\\{8y82EwbSOw>/bT9g,EM)3cyavRq8"));
$write("%s",("dEc1:ZZ>Xxly42qwZ3gWc3Q\\\\{bGw@X2*yEnv46b:Da.z==xw2\\\\}<3p4=a/yhbhbXueQqz87zEOQmvabo5v6<ak|by7\\\\{<ak|g5zP9w72ebXauw01Y2Oa@a|1iJ;xa>w|95Dam7jx/bpIBy5.gaqUXXWD33\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'3at9gbOayv?TcxxRb-jb7bWaN4Nv0MG:fRgbnvT8b-jb.wl5-3[-3\\\\{6jDawbPPk>xb+VE6Bx@MSy0\\\\}BZc1:ZEao.5H7WcNqQy8|0T-r0l-uwAQPazbRaU\\\\}NML|evnw@FQPb-Jv|0zbZ;.DNv4b1vtzQIeCUG4b1vj|DaW,5b8\\\\{0R3bW3fbuRK-t<fOAa//\\\\}bbvg,EML-Mva-LS+V+wPx5bNaeF7/qLqwZa3yTXE63-XRIP\\\\{yvRqQPDPx|:j;|W3|vdFO/6Iu0RdYO*abP,c1:Z0bg|\\\\{>1RwUExxOh.Z@yye??,zbVbYzaYL*jbVRS|o:BTy>NM,?\\\\}5oxrLp|j12H/UMQ8zlb:H\\\\{yWa*/hbW3,xa|wCLPlYW8/bl/AaTwp.0>6bH*cSxR55y>0\\\\}AHc1:ZdbVzLP,P12xRQ3qYEP@@K\\\\{qQNF.C+bq;rSj1f?t.2y55d*kJEv?5|b?Bbbeb>vGaUycLj>|B.wqQ+M+>5PdBW24LH>HU7Zp|||7wAaZagC*:\\\\}b*b7ZK4Q0oyMRX\\\\}azg,EMBT,,nvlvjvhv|Ymb6b|UdHYwr,T/\\\\}"));
$write("%s",("2N+EGkxbQXX.NJFs2@@r.eFH0GawUqOIUBVk4ry0.V*e|ywhR?/4MUakQ2,a0x\\\\}O;p.kxj04vn4Ntn4NtB+JbRa*5\\\\{0d5Pa00o:f+<Babl/c.,.3bbvxWlbEa8bTeEaP+XvOa\\\\}\\\\}o2L+jv*8@@Z3NWCQ8PX44xUblQ2bUa:=LzjXAa/y\\\\{bDaXZDaLu?a/b4Y8blzPa1b2bn.Va=aRyR4nJw8r1f+=\\\\{XXJ=*ZcSP6wb\\\\}4-R+RY1LP,PT9o,5PZMY9RJMw18+>bUKPFO/62zf0t<0R@3kzvv\\\\}\\\\}o273=2+Wt9X|UBFxa|U3UaYaHy39r20v-R+R\\\\}!![2iba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"o3j[2|pa\\\\})3(f\\\\{#(tnirP;)R3FcbF,?mI@zNaeFs6C@r0F=c1:ZH>HUHu3bb*/bNa|U<UwYxR7bTa/|\\\\{bo>nXGawUBTXFxQQ93bOaS9?\\\\{\\\\}Ze\\\\{8\\\\{*7k+5vK5aca55m=aJbF=H>hUB<||c=xb.bj=n7a5ZJ\\\\}v?x7I|*Zar2f,@a13UabztJ/bbvf6*.E60UD</b@aPambYuj.VaUx8bfN>C|84.c1:ZVajbm.<aG5Tv*PS|Yawb"));
$write("%s",(".T;5;JEv0WVA/<7-w0@ao-RaRaWaQ*hb7b+<aww4BaMCT4aAcFa5b@@2C@A+R.\\\\}YzaY+M7Z\\\\{yVzHV;Uvw/bAa6\\\\}i>COz><a+bSwzbRa.Ci>COYJ5b4vg,EMS|8zfNFanV\\\\}Z|v3-XRsCwb-\\\\}c1:ZODk|1=x91vL78Jr7;W9W<5czh.nJXao:S|XVIYzx;IWRIUBV?vf?t.5-8JvbUu8PLwGM*bkbbbybzb?+r1bNbU?D2zFa3bDa?aJ*<a5zpWHz.bX>Oaxb=RERNaX5bU?DJFo,bU?Dm5a#aJ8LCc1:Zj>S|6vPPz>QPeXRFPPz>H\\\\{53a&arx.SDa;5AU\\\\{5TVvEh.JwFHqw|Um-kC<1<b4b\\\\{a14aCuyGad8\\\\{bWK9E48hzB+DaRYN4a0bp0FMoxnYBaNa*bDaeXRFU\\\\{WZEKCKW/.9ZaXa:v*zc1:Z\\\\{C<FDaRYp:B8mIMM*z,Y<2,R|;yX3WSRM2HEKbK\\\\{a4Y3W39b1vQ+Ovz8+V\\\\}wBH5vPNaY/;VzW0KPFOE6@atbFa0DakcUb/6GP=?rvw|W/Y.<a=-tb+Dm/rYc1:Z.bFO/6fN/6GPMN6/Avd/sXL\\\\{eb5AyXwb65PDQdo\\\\}ExY.>;5-lbjCSvQvyybx3bgRcMl,tb,Og,EMW28\\\\}.bZ.C@SF\\\\}80b?06r6.f:+z5zQx;E4bBy?0/bwT00C85AyXc1:Zg<jRJ+C@SFQxtJ*b<atWr2n4apb65PDzbD\\\\}4b+VD"));
$write("%s",("5zb3U3bVH/b.b\\\\{88;/1kXebt*?0Y+1@|IU2Y|:0yXJYRVN.30P\\\\{-,w7xK-ZUa.yhbkbaClb;53xUaD|ibevFMoxpZY3c/aiJfb+H0WoxXa:E;dyT:-eRQdXN\\\\}vl,2\\\\{\\\\{@c1:ZEIIYl6cAaib-,C@|0CzBaqV6b>-B/hR46eb9\\\\}r1H*cSP6?\\\\}Hyx.X,qzU,,\\\\{5G.YAaRy:8T4aubFaDCg-?XPGP,9\\\\}DW?af\\\\}00e\\\\{Waw.bzqQ1bhb0WFMox=\\\\{XX6+G1-x.\\\\}y-77-x,=Paxb/bALT59-*bRaRy2b@En\\\\}-,uBIYTVc<x|<Z3+3xbSh@4d/aRGWa1RUy11AHkvy6<ajAjb+bHuNaS|Ya1bhbs*/\"\"),\"& VbLf &\"(\"\"b\\\\{b,4aPdUaI<\\\\{bj=hbTV?+ib.btb0R3=bHNa|UdZ\\\\{bg-/bib\\\\{5c1:Z\\\\}D?+mbp*-bn*Za7bhb1bER@5L72bBaKX|8fb6=v-FMd,uYv*hb1b2ySPL7zb*:6b*Ms97WlQzbL\\\\{|G?agb;CyXyXby,wz:0b;A65PDhzYayb\\\\{bd|r2*:-be-2+l9f68H3SrJ8PlbtJldjbGaUyhbV|O@c1:ZAwxXEcbb6b\\\\{b@-6=Vyd\\\\{*:/YpQ6rMXj1@IuDt<o7xbEcbbO@by1be24@E+WaX=+VpQCSxR4.w<h.g,EMw4>O.Ti-LY.bev9b>-cz8HV3\\\\{bZ|\\\\{vPSyXyXWwubSu=w2y,=Pa/"));
$write("%s",("b.Z(:aQawbgWsW2b|d6b*Mc1:ZE-Tejz>|SaezUayT=aC>AXczFHIUiME-PPk>1y*\\\\{140YFH\\\\}bvbjb;AvA<2i3bzaba|.w,v-R+R?\\\\}\\\\{yM?.w/\\\\}CP|Y\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'McnbevFMd,s|E6lbD\\\\}r1F>Paxb?yKLeX<=c1:ZCa8zq857yX@;7Zs-,v6UrAWHq=3bD7QaSa/b?Iux;I,Wy;JYh7P=<B8BX.-,IUpZCPUQcyaX\\\\}.\\\\}/6GP:RuPfYfBc1:Zl\\\\{T-@@aOa>PsC2KRVN,@PuC+P0Rrxj;|WvY:\\\\}2y;R+bzv/|?\\\\{XRIP-NIUpZ-bVa4;H|wFRa@3rw3xUa2U+VNHa7aB=QMVzHy8<9be|mvN8c1:Z,15\\\\{?XL1aYoCORo,5P5URauDr1Y1tBaAaqwPP5\\\\{/z-zQMqB7-PS5b,ZX/VaTAaLW4TaLAHV;U<5Aa3be+6UrApAe0uUiBj6a3am|7-+Uc1:Z\\\\{;HBa=-AXbRae0COMU4;DaW75||BVGRae0eXzFakaWLDaeX2|Nt.FbpaB*0.bOzf+2xf+o,LNama2C;BLSyBqAn-)MAka721(f\\\\{#,43zNBya201(f\\\\{#(ntnirpn\\\\})215(f\\\\{##OBT4S7aW73=Wa7b.bRay+,YgP\\\\{,;vc1:ZjbGAa=PA3bt2@a3bz.q??af++Saea*b+>HJaba6S7d;a3bYHuGe-WaWHTAh0lbv0lbGA;BlekR=a>v<B+BT"));
$write("%s",("afHSa7-WaXA3be+BPeoavY:-8<WaWaW-jCiIa)cK-CUc00>yX*J1*BYxR\\\\}FC@@I4;Dadhc=x>*.y@DPXvROy:xSW;R9WaxR55GZxYp:vdFOoYe?\\\\{-vd>PpYtPHUPNaYivVzc1:ZL,qYVOzFn-vdFO2CwYo:|BP4>TwZ,Yyw*b\\\\}59bzbEV7-d<RVTahc-\\\\}4;fLvd>PtOfYGVc=oCmZ?J1b>K-byye?d|/be|Nw\\\\{KRVwz0yaCo-c1:Zles-z@a?a:\\\\}2y55iPkxfzW;RaWaWa5wvySah=WafF+bWA-cWa2URaWag-SaVafF95OS#3e,ZaMa:z9\\\\}/b@5k6p:M@4vOa/bDa;5wb,9lekbk<6b+bIFoNhJr1CS4xCS0AH>eYEVWaOaWa2U6bd4Q3aYe5v:+oR=\\\\{|CmTRa;5wbh.YaNUn=UaB<SJd=iH,RaUzWPau*AZT<a|wek|uz1baCvb2ATExHRIrwp-g/|,R.A-7N;xbF5OL\\\\{++V|RI1bI2BEyb6J\\\\}b5wE6-0P01bF0Y+E2R5RaW8hR46swP6S|y*wb@w6b=a-U0v6Ui4iJ0HkCUa@aH*c1:Z@JVO|1.Y5APa\\\\{b*V+d78<KW75|+F<MzRf:b\\\\{?+=.5xUaU,NaibfZ++leVaJ6zBI/3\\\\}|Lmb|ya\\\\{CKAaEDH*cSxRrx+wC=o|ezUa0HS|e\\\\{l7+b\\\\{bPGEv*P3b\\\\{8TL:CEwzW;3ExuGS|j.hb\\\\{8F<P:WyD|\\\\{b"));
$write("%s",("K5VbFayb2b*:h?-2kvdbeTZSc1:ZFcUadbfH1bqw<ag3,b@+Far2t8j\\\\}EI?+?x;5G.t<AL\\\\{@@xX47=7ySu8JybhbmQiVYa0Hb*5bbC,Vcwa5HR\\\\{yT:-aCCYSvgP\\\\{,ePlAXLa#a3b*:R7?+0b4y.SYuFaybzbUx\\\\{Lx;?v75apbl4Fvt9FctJfH@6E/r1o5c1:Z4A.wuvz5K9L\\\\{C.mQ\\\\}bDarzjbS|c9QRP,9\\\\}eb=aTapQ+bTaFvzbxy>ZYa|by:s9T>SR<aw66b@a9\\\\}+z=3acbYaRHs*2.6FK9|d6b+b3|bzHR4b@5lHdd,,8HU.M+3b>;LSzx;I=PB8PNaY,?uPfYg252aUdbu?s?5*V2@U\\\\}8c1:ZDXABla(f\\\\{#(tnirP;ECBka3(f\\\\{#\\\\}i-zT;Wardu@XIRuPuvdFOmOG>RybbO\\\\{wPA.3bSa/\\\\}qQ\\\\{yVz3:Vz5vRWkCe.t9,b=RTY2b?a|z.bGvvBhbUaY52z>C;7HVe?zE4ZCOVOr7;W.7YyDaNvG<Cwdwmvk*0TqAtJcb:0R4nJh|NUf>QWmv=ac1:Z+b2GSaCadvt/LDmH?aSax|M@ayfb?|g33bab;J+bB\\\\}fH1byDSG7bu\\\\{le9buy2y.b-V7bs<X/tscb:3d/:zv4-<ubSaCaWaR+t?-4\\\\{+@aabiR1*lbq8gC+b8V9b<albbbOD*,O3gsae<;xc51<+b2GW.ZU5UJ4a\\\\}aq8y6y|CBjRwbd/5bhz"));
$write("%s",("1<+bKw:8/5o3apbC*+bk-|bs<Sa=\\\\{XX*IE9H|X3p40Uf/7?CaX4|4ZTS>Y.:0I8nJP15vF?vbYGzFCa:><zPBp:SWe.4vbb\\\\{bZaUx8b2b=EkHvwyb\\\\{btb?Aa,bDa/1L-Mv|*Za7bzbF?eb4EGa<H<ajAV:bbe0RYFHawCOe*L||U<U?ziH,Rc1:ZAzI|0b\\\\}wY+@.D*lb14o::-C9g5+>5PGXE\\\\{3b3b;?UxYUpO7=cM7-z@v9e0RYp:GH)3aQa*z,Yx;QLDaNv<zCa|;Gy,wAveXVRaz\\\\}:PPz>IUpZlGf\\\\{F=H>hUc1:ZeXn>|WaIp:kDD\\\\}JYleV<DaTNcead?QPk3cRd*z,Yyw4@j,TQS|rYE\\\\}U-s+cSRvEaCOiYHVe?WaXJyy4EO-Y=hvc1:ZkvFaiCK-jb7bx|Ca\\\\{bg-k;K2/UK2kbFavfTaxR<.iAS\\\\}Da/1d04:VBP614/|l7K2-bGar*p*-b=aC>1KD\\\\}5vVz7\\\\}.Zlb@6jvS4m5yXwb>-TW;dL7>-tQ?a:7,SW\\\\{=albe\\\\{O2TYSB4xV?7NgWw;,x==gKCaz8\\\\{-w|A8kv|Ic1:Zxbhb;E>wBQK8Gv;E3Q,x4@0H@+GKiKGv;EYAw5tbDND6>a5-Lztv3\\\\}a9EauDpJ:Ma>h+DNIUD=9-fb*No.5Hm53Wl*8<IUBV0WFMd,|-TAh0\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'tnirp*P[4@2ya8361(f\\\\{# wohsn\\\\})2575(f"));
$write("%s",("\\\\{#0B[R35da442E4E>6Tka;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\})00611<6[R39ea0603F4[R38(a93332(f\\\\{#\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\',\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(rt.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'jbYaIUD=o?OX-XWw#@auc65leY\\\\{W\\\\{U,F=H>eYSF2bm5JYc1:ZC9wbe-v*\\\\}@d|yb9V7V=V+VSaLDFR/b;72bw-Q+nzPa/bhbW3I6N2BaPa?xW3Va\\\\}df/@Fe0B<*ZcSxR7bTamv=a*:*FrwL|\\\\}57|W3ab3brz\\\\}b*b,.IUD=AT4b@*,Y<2Wwo,5PFT*2leY\\\\{0R8\\\\{2C@Ac1:Z+R\\\\}FqYhBaYqYz>DWc2bZNrwBPVzLPlY|X9bhb,bTa|bWwg,EMA|+M\\\\}55vzAhbvRqQhv|Ys-2\\\\}nv-e;=xwvw2.F9IY=\\\\{XXmRIYTV4\\\\}NuSwRI2Qlzq|OaX\\\\{d8Lwb8Z7ebL-L730w6pQcbe-R?z+t/jO|>3Za/aOx/SW7NKC@TR1U\\\\}vKQebS/dG=a|UdZEaRv18n.:@2b+3c7aBaOa1U\\\\}v4:9V+Q4MPRSES9Aa|UdZ\\\\}dN@9V+Q=/C@fw1UTuc1:ZW3cUe-wG@mbV22:IYTVIY/JlC>a3Sjv+Q4Mm3cw7=O7gbl9kEXTjEN.jDjb+dlDf:dLTA*F3|Pa\\\\{bmI@z|YPa\\\\{b<RqQ\\\\{yX\\\\}wbOVud0v6U-?q=xOh."));
$write("%s",("Z@:-N+L\\\\{G.yb+Vc1:Z6Zd/:8zW5I7bX3nZSEZ|7--b<FsBsLO9|d65/0cZ,:zYS|6ZBaGaKZE\\\\}*.bv6.6QTVIYTVRW1vlH.Zy=sLW6\\\\{b,S+e+b7\\\\{vbAYHu<ZuT4bw4Yy6MQMr0=E/U1*Uac/h.3,w4E6ibr/GYr|BYYaQMp<EaK-y.jAKb0T-b2bYam,H*vZU7fHN0LJ.2y+bXbb:8sFw0HVrKzwiL-W\\\\}L6=CM2KeyfvT\\\\{eH2bY+*0ZaTR.b@akbI2|S8b0\\\\}n4?\\\\};\\\\}WK3ba/FvsB,U\\\\{X--uXsB?eVNxS+V43s*m2G0uR6ysXOz1yBa+yq?[R39Z0hR4EEaUaN-SG.bS|xRz<6RnDtR:z3|Cz5|l9j9-wy>I-N+4wubJPnOsOR3@PFP/w@32\\\\{oOA1ONrO-|c;mOsPf?=ybVAA14x9e|j.?\\\\}l@n5zK\\\\}5:zf\\\\{9b2bP1.QU5Za6WS4.CD>GRGD.bCaE2VyQWUMO/8yd@7bOz2vj*Hvy*h>xHI7a*lbEwiCCaC9zXlRSVybWw:+VV-C@aw8\\\\{1l/cbG18zAa6y-b7*3wA|DOmV4zz<Z?z,?Wt-s.ubLwgb,be|x9Raw.pW,.Gvs*O.*v|12bUSEa70+bf,I6A;60A.Ru-,?MjbWa|7Za>aEaz|oFnHY2@5cbry>J>xOP6b<.hSlSsG.bQ;XyVyBP?aOaybYuD5vb3H6bTa@xg18zk<Avkb4x.wa;m*lb6xczb*=7Q\\\\}p"));
$write("%s",("Uz@-UPSmB-\\\\{C8fb|EK\\\\}7*sSr,\\\\}wCVGBjbRa|wjM|9eVa>=,QuLS4vO;Vatbfb\\\\{Dn-LvYvAeF6m2?+QM-bQa5vTaiPJ6>@ByoS0\\\\}j,QUl4T||8:vzSkNr7U-3-vSUa:8xb@albt;Lzz,W.YP\\\\}CG;1x9?NE\\\\}bib6yn?YwCzUSEx9F\\\\{>qB\\\\}</<jbiU\\\\}G,.aS>wS;Ov/>7b6y4bebVyf?B|WauIx8/vGT8R4vNazbhb?aleG9EI+U7NRw,RGa1fHvjS=Hr1*/RaPaK2Da=\\\\{pTsAeI6y3KaB5>aORKj=HIbLx8d+tM4PU>Kz\\\\}v,66y4/xPW2>5A|x8USfNXvsT9RT+?T71aN=T\\\\{>j11<kbYarSmbLC-2Vbe>sT6Q*yjS,E+z;5iLmCe>Na+S-:n?O|7*@Mzb-:4;QawbByy*/<ledJUS00=yfSe\\\\{\\\\}z\\\\}bNa*d7=,.t\\\\}YvcbOaCvTSxv2*Qa1bA|6bgx\\\\{|Y+c/=awEOSkR4;GaNPA|cf,.4bJ6N.,SOMCa90A|\\\\{bdb-|LzQaizv92vg-hc*dY*fblb;1OxDaOz6blbBacNOziz;E2vzwdyfzs+CD@:wD*b2bAaNakbwDM0CH=|2vs.F=YPnRc\\\\}*zXMjzA|TMs+jIlPfbt7Na2bP=cbiL=J@M3b6wPa=aAa:>0PPa2bhbuby>>KAILBvbTaTPc=vvmIlHJL2RTxUMh>JMGa,zSP/vAD?asM@EX.iv6w:M?\\\\}"));
$write("%s",("ebIxnDWaIN:.=-M@Q\\\\}aQYP<71PYGzb+bXaT>UN7b=aB?3b@-*@x/2b4QlE\\\\{v:M/bPu++FQOaDQu\\\\{wyf+Oa7-fQf+x\\\\}lzo;A-\\\\{\\\\}ub?w8QwQ=?5wo\\\\}zQXy|2\\\\{v;87;Y|q8q|?.B-M|:?MA=-0bj\\\\}Jw2KcF=-D3=?e-KIv\\\\}Gv=-r,Yacbl,-bOa8bD;,xW/8-zv?/3b70d5=\\\\{*C4anPFz=-3b<A.wmbtzDaCO><wbM,\\\\{\\\\{>AuOxAKGHOWOEOkvE6dbTa-PGOV1BOf?wOuBF?|bjvd+hHID3\\\\{<8MHFER8Y1eBM3JMUOl99F@@?76|Y2Wa,bJzi2NN4-U@+K|OzOtN>8=?,.lb,yQwkKibXLPu1yIFOOs@Q3oOOwbb004=\\\\}5-cc=PLvwi,Z|hc?HEzvC*3e3wzzxtN<AG9ByA|kbhbxy|MmNcbTE12qFWa@FdA:/5AFxfOu/v\\\\}dy6.\\\\{e2J1NPa/NZxr1kJj\\\\{tCx3nKc,Dxub=AKxc3x=HLOaIF-xyyDa\\\\}bwbVyXxlLl>NK5.v\\\\}wvcxA+8@-/pKYzwxmK,6*,Q5Yadbf?WJeMMwKwIw?NX<H=I=e-?w=w-\\\\{058=:8RL9>5w3w4a,IyM@dwM7b*N0w2w,wD41@84a\\\\}W?TCe-C.3-*LUD-/+/\\\\}/CEtyry8z=6?M@yCacN,b?ECv/>X5JD\\\\}>z<ILT1J6RFH9Jb5-2b*d.v\\\\}5abH*yH:I@xNI7b+GG"));
$write("%s",("xLwwy0\\\\}Ya,bO7O@X.6Ewwxvb*O.oxv\\\\}7zXa78WyN-abv\\\\}i.A.9b*b?aywuy4BqH1Lvg/L*5iH-0gH6beFyyBv\\\\{>b7KyXxSK>IYybvfzsI;xNKubjvAH|8\\\\{\\\\}zAMuHy+d5:\\\\{K+vRaZ*25+\\\\}h|\\\\}4\\\\{/g>29;=/K6/f?wLe7bbwb4.7=7b\\\\{+.|rIZJv:-b7bu|F=.-oG,Kng*KV6??s2s+@J|3,b+d/>DKh7qCi9675ItbXa0/hIbbA|e\\\\}i;U6=,PxNxiIIB*bZa?aSAEaPIlb00cb364DX6m>Z5/1y|y7Da*@39zF6\\\\}m7.xx\\\\}W4DG0bBGXbhGYF>/\\\\{,kvfwhcrwNj39PvfwK4f@=aN?C2X+K@4akF3J>f1J6/3:wEXG3yaH,c83V8G0f?b\\\\}+5c;JxgB1C|,z,LwRa.b=adG93T\\\\{a>rIyb\\\\{>zCr1-/|6X.+|NaEaVa;<mb9<|wlJ<J:8Raf+i1g6=?;J2bGIDDy<1-TET9VaRaH6WvOwfHh|nFYD-IKf+Im?lG//*ycf\\\\}b+b|IWvK8vb/<P6a\\\\}pv-HNa2,jb4x3bQ;X2\\\\}.@B1D+H>aQaibS5F0NajxK7j5i+VuTuK4s.S*Wac/VaBa4AO*v-I|yvY4Rv2bRaTA:8LDv-k\\\\}qEx,Vaf?v3,:3-=DW@*.X3j9@5ZaMz3/V7X2s.4aeDrH-fpH2bx,ab1\\\\}mbu\\\\}30A?7|@a.GYv3?2,Aa:7X>LC0C*z"));
$write("%s",("X@x<X?WvU:/z7vg8-b@xSvNAr6Va,.m|-bOxdb;5|bibCwvB07c*6\\\\}Q>f\\\\}\\\\{b.CjbR=G>Z.5bBxmvO*le|bO*gbFc1bT+Z-|b4vc;@aRy+b@5YE>ay=.b=|Ev1bg|@*U9<DB8-4:wU@1BpGffnGA=BBfbzb\\\\{>e+*?@D23lb2\\\\{\\\\{y3y3bJ23:6FL@IGXbebm7d/eb65Zat-r-gvw@eby:;<yy5?w\\\\}p.mbXu0bnEt@gGS72F0F@\\\\{nzP+WBKEs00.>?u8Qvf:7|||d;evvvf,h2J1lbu\\\\}.7q|W,E?39UaF>N@S<CAlFrejF>aWB\\\\}/9=Tu8Fsv2\\\\}a-ewY5f64@kE4FWwfwvfVy|:Ya5bNtWawbzbkb;</bubLCP3v-e@lepy\\\\}vvB9s|4Wv0?W,vbNDnEwblED>gEsv-,R7x|jbp3W7k:i:OeED/bU:O*s7SaZ7t\\\\}==*0J?C=6ba50ba>Bw4aR@ZDfeXD9sLCr4Aa\\\\{|U,e0yv6xZ|qAk9TaR*,,7Dv\\\\{TuvfcfGy-,-bExj,WyGaZ\\\\{\\\\}DTa0E\\\\}\\\\}.b?5O69-Ev-bZaJ5bb5bhb3/jv7wN9kbdxJ*H6+\\\\}37p2mblejbu;|b6b0bbbmbo5CBpvV?T?6\\\\}p758OCP\\\\{TuVu\\\\}v.b<.T*5A;CSam+-ba>s/o@fDSgdDkb@3Y?s6r7b<p37b@a;@wB\\\\}Dw>.Bw?>xyb4vew*z\\\\{C71W51x-BH*Y8U1P4-5K>Qxn"));
$write("%s",("C=*JBa\\\\}h7w-Ya=@fwaw@-y:v\\\\}NuRCJ?Oak0=aibo>-bNa@aj>E/C/S/\\\\{+wb30ub+bK-Xx4az?2BEg0Bu.Y+C.DaD7|bQdn4V?@\\\\}o5:Cl/g+b-rC\\\\}4sAe2w\\\\}@8o-Y2zvWu\\\\{b-86==;ebK-ybs0?=9CuBXB+6A.A+F984Zz*=.6bbaz|4\\\\{b@*=yVt=yh8bBXa2/C8Y1|=W1I,+4\\\\{b+||b-wOxB1/3,bYy*bx|=aM+aw-y5vYv,bLw\\\\{;4AhxYaWagcYac5wwR.S.Qal6-b@36,U,f?I\\\\}-53567\\\\{@x@>\\\\}9B/bh@LAr1P|j;/AQ*bbf+/v4a=>DAShBAU=33r>OaQ*?a3bU:B*9=U:G<\\\\{5sBtBz@zAA-Sa8bnA97K?v8I<Q+@3L1b3\\\\}=?Av/N8p>Ga\\\\},Wa@aVa3b2xfbhbSaQ*>aZ:s>5@W4jd9\\\\}y.W4f?4aL=S@IhQ@5b|\\\\{o132\\\\}3Axxb1v1@@a8<=aM?O@TaebQ*F=bAl/=af+Q+a06vA-p?N@\\\\{>,w,c,bfzt4.?Rx2bR+t-=-0/o:6zXan8g.9br,2?M\\\\{o9Q!![2iba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"o3j[2|pa\\"));
$write("%s",("\\})3(f\\\\{#(tnirP;)R3FZ0=cxbbz<z/L8L<4aP<p@vhn@?=y@M@|@zbR6;8g5ab4b6bXa|x=av7t<,bYavb@aTap4f:0/b\\\\{l7|65.Xaey1.A+I:U,MzX75wU7=af<o?O?L?M?>=eblxS0wwR8O=I;\\\\{?>gy?Z==aR+Q5nz8b<.7=4+j9U,cbN8o6:/U,|1CaXaOeO+*x,:T<N?p?:>n?,bWuy|MvI-absvB,0\\\\}<656f?g7J>mbkxY:o1W:ayleDaibX+/.cb*//3V=*>U.Wa\\\\{*U=4a;:>>ph<>V5-6?yT\\\\{3bYwi,M<D>?=m?C>b;0\\\\{0bh+S|\\\\}w4>gvc=y.b;Lr,.tdjbB+lb\\\\}v,bnvQ+W|8zyyT1Y+0.4,|6M0y=x4CaBwB>A=A>L<v589M=RgK=:8B=/bTz+e><|w@<*5o;Wa8x\\\\{bVaR14vo,v>s9DaA0o>r1fvd+T=b=W.X:j>h>T9Yas\\\\{E=?<U:fbEap612Namb2byv60Ba<6jv=,bv71V*V5Rzz=x=mb4aj\"\"),\"& VbLf &\"(\"\"8Q<khO<gb8bf+N0b6n9c:z;@=U<M<V<FwdbsvOwkb2b@-ib/b|d\\\\{yUay-e/Rap5m|7<.bJzS3q1N3\\\\{4W6vbh;1zn7r-EaabWaTa@aW/SaTaWaAaSaAaOahzTa=amb|4r1n*VaX/n-4:h<T<f<4a86J;MgH;?9|;g<SaEa/b;<=aEa6wQa95VaXxd:?8n-Pa4<Uax8WaEaSaW4"));
$write("%s",("2y/<Val7=aOdTaBamb@aWaPaWad4:5V9M8@0.b9xp4lbub29q8y*ozP;n.Z+Yv,5B9z;e<x;d<\\\\{;98.bN,tbN/lb\\\\}5w7+e7;wybxdbK4mbewg;4as5<:Di::hb8xVutb/+Z6bbibEatbB/|+z+7bC32b1bSalbk*eyn3Rag;dbZ*-.s9mbb-z5y;G95:w;3:D9-vF-r1\\\\{9X|l/gb+bS9o-/+p:s\\\\{y4m9m:ZaZ*Oa,bcbNjP1L|4229Nt|4<a8\\\\{Y.nv?74.2|7bG:.b-+Nw2*Ya=.K8r1O4-9cxtb9x;+H399wi792/j5=aD94:H92:F9\\\\}5i-x:t\\\\}eb5b*.Xa|be/e\\\\{\\\\{bmbjzNtTaP2F2W7V/\\\\{b/0r1l9Su+\\\\{B+SayvOa3bk9e\\\\}\\\\}9i9@aNaB-Pu<aZvL.R-X8ew3bD\\\\}?6VuRvtwv-Eal9B9;8E9B9?9C9:8=7>9o5<8Sux5T8>yw2k8sji8cb?aW/fbibA8TaO4ibVaYaVas\\\\{a6Mz6/y.,.+bHvZaTvF4tb=aVaFaM0V6E.BaZar1=a.bZa18Xugbs-db<a*zK.y/B/AaYwcxK-kbXbabe0\\\\{/,1k1Rakbf+o+7brxm2Yw-b+bRvr1@36\\\\}z5Aw:7;787\\\\{,.bebkb|zuyY.abjx7bSyDat\\\\}F-4blb>aeb|bmblbPa8bs0NwD.A/BaQ/84\\\\{b4aa196mj76,bRaFxEw\\\\{bM+V\\\\{1bVa\\\\{7f0Sajx\\\\}"));
$write("%s",("bbx90mbC3SaZ|5.jxzbL-R.14,x0\\\\}o+OvVa5.Z|F\\\\}6yvb05<7n5679705Va>a57z5X,fbz5f|Hukv1bh+wb?5lbUuhv4/cb2/pvw-QaO*XaxvUuY2j\\\\}Qamb3bF4c7a7Y6r1ozE--.:v3\\\\}cb60,bDae\\\\}G.h2K0Yyr,..V|-b\\\\{bub;5ebY/>aibR,X,Fawbvbg-Zaw\\\\}u\\\\}k+ozx|*b4ap/t5Vir5/bjxvb;/5,mzKzw3Q3vbhb@a0.+525Ev=|zbl|Oa+bE5\\\\}*\\\\}52bzx-1B1\\\\}w/b?5kbl4*.@a=-ybvbf\\\\{|wz4L0@\\\\{kbo,4342J|@aXac/Dar06yUa8-|*v*a/j,;dOaB-f\\\\{0bDak|:.kbPa4b?/UaEaEaAag0\\\\{b/bWas,q,\\\\}5Nu\\\\{5vbAayw*yfz7/|4AwBwm5A+XaDa4a+-I3|iG3Na=a>aGwCwgbS.RaB\\\\{ewlbBxgcyvVa7*ZalbAalbgbM/K/m+wbf+.v3byv4\\\\}O+mbOa3.6-\\\\}bkxO1JzAaL+LwWah1Kw=a3bLuWw3+0/:/oz8|U+W\\\\}.2weYaP*k1Tafb@3Q\\\\{azDas4Xx=\\\\}<+a3UafbFx\\\\{*61,\\\\{\\\\}v\\\\{b30tb+b>aTa0/g|r,RaVatsSa?aozNa,bhbCaZa6b2bf1K1Fzf2,3m\\\\{42N1bv4a8+x2Liv2U1vbs0C.*+u*A0;*O-k*XaXwwb?acbm2ubd+x*o1U0Va\\\\}/f|g3\\\\}b"));
$write("%s",("dbf2j\\\\{y3NvE1x\\\\{l1d3e16ro+|+\\\\{y*+kv@-kvn.4b*b0bc2+bkbQax\\\\{M1Jz@1h2>1iv\\\\}bab0b=,\\\\}y;,G1UaUaibUaf/0bD|lb3y+b6b,babwvfxZu,b=wB\\\\{swswGal\\\\}Fw8\\\\}SaNvvbY1p1V0K,C1J.wzrvfb4bn0T\\\\{/bBafb:.4aO\\\\}b1@iZ01bUayblb\\\\}\\\\}vb?aBcibg\\\\}u1f1Hxnxn\\\\{X1.bI12bn*Y/ebVzL,x\\\\{h\\\\{+1tbjvYykxgbV.m1B1Yz?15+8xx1>aL+M+j\\\\{w\\\\{7,JxHzd,;\\\\}gz*bmbNv:.e+7wn,kvRvXyV/mbCaMv?\\\\{G*=*w+EaU,\\\\{b*bfw2b7bHu8b6bUaN0<0X0TzTxy\\\\{J,v\\\\{CaNa|b@a-bJxXz4a;\\\\{q/Cio/ebDzBzz\\\\{v*YuWulzwyab-,jb/-F..*UaFx>acb\\\\{bibxz6bzx2-rzlbU,|w|.Aal/kbe-z,Aaqze0n.BawbUaFaTyUx8y1*7b?ePa.bF+D+0bUa5.R+5.BalevfevS\\\\{ubP*j\\\\}Sa4bhbWaUa8bEab-UawbkbVaSa3bYaQv3\\\\}o+/b/yNyu,l/ibdbXa>ve-,xmb\\\\{+nw?+TaH+mb+bb-lb7bfwA+//AaO*V+jbXaMzWau-ww+v@+Xaa\\\\{nzcbab/bfbi*9,F*H,+wB\\\\{m,+bx|4a;y,-/i*-ibTwgblejv,\\\\}x,Oax-XaQa4bvbUaZa8b3bM|K"));
$write("%s",("|-bSamv*bS|,,A|8b?\\\\{r+8,E*Xas\\\\{q\\\\{d,lxNvibLwdb1\\\\}-,FaOa1bm,/b6\\\\}5bO\\\\{8bOa0b5\\\\}=aOws,+|FxTaFar\\\\{0b>+u.e-8-AaUalee\\\\}/*++Par\\\\{v\\\\}lb0\\\\}cbybNaUx*bibjbQaWvtb,,ab|d\\\\{wfwQjr-5v8wzbdbk|>*Ywt\\\\}x|/bEaXaZaNj>aMvj\\\\}Ua5byt|z2bCadbezkbgb*b\\\\{b?aNa8b=a9\\\\}wbDatx/,-,|w=+4alw9+gk7+NzWaXaOa2b=atbcb8bwb.bVa\\\\}bSauble.bkxTavbvbWaQa-cCaY|kxebtbyyQ,*\\\\}Xapzp\\\\}DayyEacbSah|ZyDzl\\\\{vdi\\\\{=*.,**db1bB+lzu\\\\}zvuwOa8x|bN*Va?\\\\{g*\\\\{zg\\\\{b\\\\{ozabcbAaj*s+x+ubgb|bnzle8b+dbbkbWa0bb\\\\{bvV+X+zbWaV+0vW*c+8bmb\\\\}vzb=a6\\\\}IzPavbo\\\\{Fxvwlbib>ayw>xFx.x*bzvRa8brvabRu\\\\{+2bWav\\\\}S*Q*svRvxbEaXuvbVa,bPaXxd\\\\}p\\\\{4aiwP\\\\}ckN\\\\}mx+b0beb\\\\}bEav\\\\}ubAa>aqw/bv\\\\}zyBaeb8b*zq+D*BaA|I|h*8\\\\{f*Pu\\\\}b3bZ|NjRvNjXukb3bubDaz*U*@y@a\\\\{|az/v-wy*w*TaAambgb\\\\{bAaivub7biv*bEah*?*>x<*Qa@aA|Avyx7\\\\{hbzz"));
$write("%s",("u\\\\{XwVwYa3bTaQv7b8x7z0bRas\\\\{<\\\\}KvRa5bo|4b\\\\{bjb/vPx-b@aSz7bEa-blembwbvw0\\\\{jbEa2v/bg|zx/|\\\\}z6\\\\{f\\\\{ib\\\\{bAx\\\\}bzbTaXvSakb4za\\\\}+v4aXt<\\\\{Ek:\\\\{6b>aD\\\\{C|wb2\\\\{ib+b,bdbX|V|Xa\\\\{b7ve\\\\}r\\\\{c\\\\}/b1bPa*bNtcb,bWaCa\\\\{yEa1bK\\\\{/bdbcbWa.bg|IyGyrwZa/btbgb.bAaVzPaa\\\\}Da8bhbVy\\\\}bmbBaXwrvQajbmyPzNz\\\\{b1bdb8b.bTaQaOa\\\\{bUa+wab>a\\\\{|kx4xhbSzybDa.bqw3\\\\{,eC\\\\{A\\\\{Satx9b.b?aebS\\\\{kz=zVa5bRatbw|-w!![2iba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"o3j[2|pa\\\\})3(f\\\\{#(tnirP;)R3FZ0YatbRatx7bR\\\\{\\\\{|ozSaWvAaEadbSaBacbmbmbXa@zrxcb\\\\}b.b,w/bVakbNaxbYufbkb*bTaNa5bB\\\\{levb.zGa1\\\\{mbevzbNaCaNw3bPuxw0bPa.wNvybRarwCzOwle3b,bhvEatx4aTt<y=k:yvv,b|zv\\\\{xz,\\\\{Cale-b3bU"));
$write("%s",("aGa;wRa0b2yebm\\\\{1x/xk\\\\{9z?xMxYa\\\\}wQzNaOzox*dWzUzSzubBx@x>xyzFaebOarzmb\\\\{bKzIzGzEzgbCz?aAz|wWx;dNaGxib,bEa7bIxOaGxebTa4xRaUxjy5blzjzhzSa5b.bAx|b7b-bFa>a+bjbUavbzblbleebEayxGv+bbv:vLxQazbWwRazb=wXaSa\\\\{bWaVaFxubQa\\\\{b.bUaab5b<aRy|b\\\\{bkbdbvbOatble*b@aUaQaPayywyhb>a,xoy>wNv/b=a1bRw7y5y-bFvdb0b4aPrjwukkwRwib0bZa\\\\{xUaPa7bDa@aFa1bWaYvzbAatbebmbibTadbmb.b-bdblb\\\\{w,xabyv|w5x3x1xSxTvjxbyfx,bdxOu*bXaEajb6x4x2xFa0x.x|b/bAx2bbv=x1bEavv>apxvxOaYaEavdYaFa.bhb?v9vqv3bAa0bdb|wWagbwbVa?aNwSa,bfbcbibowdxbb|bDa>asxqxoxmxZvYavvTaOavbZaBaBv3bXabbhbNaBaDawvtbabubhbTaab.bmbivBbjbPa,bAaCaFatbWaBaabwb*bqvNujbleAwDahb9wgbvbNa1ble7b<a>adb/bSaXaFagb.w/w-w+w/bYagb7bzwjb*bAaFambSaYabb,beb1bfbwbbvWuAaQrGjhwUtUjWtXacbhbRaubWuEa>aFa7bNaCvvb2bXaabzbEaCaeb-b/b-beb9v,bNa7bvbCaEa5bDajb"));
$write("%s",("abjb.bkbablbzbUagb5blbjbdv*bjbDadb+bmbDavbQdZamb=aYaab,b7bmbdb.bOaCaDa|bEaYaeb.bWatbdb5bmbjbcblbhbjbOu2b0bcbwbSa1bZa|bWaubabhb<aCabb*b7b?aQa\\\\}t4uds1uFt/ugursltVsSrJsnu3ustzu,u;aVsPsNsye/t;tJt=tpuxu-bVsutCaYsjuoubuwbWbVs,tssng0tduPahuEa@arsGtcu>tBsYsLskt@dEt:s8sQr:jSt9aQrkkOr-b4byexfubjdTrpt-t3tmt<t?t:tps9aEaOaJsvg4t+tqt5titZd:a-bJsngot=aZs>frt?sdtvtfs1sWs*sUs@a<a-bTrEsQsbtZsKfXs/sjtct\\\\{sWeysJs>fHsat:aCaYrIsDs>aAa-a-fqsKsws|s9a8a4shsus?a>ars@sZr>sKf<sbcYr=s3sFaBaWe0sxsjs-f-s*bvbtb/bye:fTr.s\\\\}stsyebsosDrmsOaTrnsvs?aAayepsTrXrgsAa@a-affcsasYrisWr9aYrHareMr8aCa@aWeyf\\\\{bvb8aSr0e8arb8a8a2b4a4afk4a4exb3bCb6byeDbbcubHaff?h-f;fAhBh.b4eQbye,bMbKbBb?aheeoShvr/rqr+r|rsr*rerbrwroruryrnrfrrrtrprmrAqdrZqarkrlrirYqjrgrhrUqWqTq=qcr7qRqSqXqQqVqOqLqMqJq8qPq5qNq0qHqIqKqG"));
$write("%s",("qDq*qFqBqEq?qCq@qvq>q;qjq:q<q3q6q9q+q2q4q1q\\\\{q/q,q.qbqrq\\\\}q-qxqzq|qpquqwqyqqqtqeqsqnqgqdqkqlqoqZpmqUpiqfqWphqIpFpaqSpYpcqRpJpVpXpTpQp+pHpDpEpOpPpMpCpNpKpLp?pAp>p\\\\{pGpup<p=pBp;p@p9p6p7p4pvp:psp8pnp2p3p5p1p.php0p,p/p\\\\}p-p*pZo|pypNoxpzpqptpwpippprpopepmpjplpFoVogpkpbpdpfpToYoapcpUoXoIoWoRoKoHoOoPoSoDoQo?oMoJoAoLo3o0oEo=oCoGo<o4o@oBo>o;oco2o.o/o9o:o7o-o8o5o6o\\\\}o+o|oYn1oSnzo\\\\{o,oyo*owotouoroTnxoQnvoLnpoqosoooloFnnojomoaokobo>nEetbLjFg:lkkZnWn2nVnXnOnRnUnGnNnPnMnCnKnHnJn*n:nEnIn@nBnDn8n=n?nAn9n<n-n;n6n/n,n3n4n7n|n5nwn1n.nyn0nknhn\\\\}nun\\\\{n+ntnlnxnznvnsnGmjnfngnqnrnonenpnmnnnancnZmCmin=mXmYmdnWmbnUmRmSmPm>mVm;mTm6mNmOmQmMmJm0mLmHmKmEmImFm|mDmAmpm@mBm9m<m?m1m8m:m7m-m5m2m4mhmxm/m3m*m,m.mvm\\\\{m\\\\}m+mwmzmkmymtmmmjmqmrmumfmsmamomlmcmnmOlLlgmYlemimXlPlbmdmZlWlBl"));
$write("%s",("NlJlKlUlVlSlIlTlQlRlElGl8lAlMlvl6l7lHl5lFl3lDl1lCl/l\\\\{l@lul=hre3e9i<gJjfl.lwl4lql2lkl0lfl,l-l*lXk+l|l\\\\}lzlNkylrlxloltlmlslilplllnlbldlaljlglclelhlZkFkTkWkYkPkSkVkIkUkRkKkHkOkDkQk9kMkJk;kLkEk1k=kBkCkGkAk>k5k<k8k@k.k?k*kvk:k/k6k3k7k0k-kek4kYj2kZjtkuk+k,k\\\\}ksk\\\\{k|kykqkzkwkxkmkoklkakrkGjpkUjnk:jjkkkhk1jikfkgkdk\\\\}jckVjbkEjXjCjWj=jFjHjAj?i|b|bvb?e.b3b>b9dJg7iIh;jDj@jBj8j>j6j?j9j-j4j<j7jtj5j0j3j,j2j\\\\{j.jyj*j/j|jljqj+jzjwjgjrjsjpjkjxjujvjojijnj5iejmjjjZiWifjcjdjhjbjYiBi3iUiViajTiQiRiXiPiMi-iSi|iKiLiOiJiNiHiEiriIi@iGiCiFi/iDiAihi.i0imiEhzbDbxfrbZdhgIgUgwi4i1i2i*i,i\\\\}ibiwi+itizi\\\\{ixiuioiyijiThvisikiqinipiliXheiiifigidiWhciZhaiPhYhVh,hRhShHhQhNhOhUhMhJhKg*hIh4hGhLh3hKh/hwh+hFh5h2hlg2b3b4b/bHekfng=f-fefJcWetf-bMgvh0h1h.hth|h-hzh\\\\}hQgIguhph\\\\{hxhyhrhnhqhCgsh>"));
$write("%s",("gohkhlh8gmhRgjhSgPgihMgKa\\\\{b;a.cwbldIaXbVbTb0a9dAgegSgNg1gOg/gLgFg+gEgJgGgHg@gBg?gDg<gAg=g4g:gwg;g7g9g-g5g2g6g0gsg|g3gxg,g\\\\}g.g\\\\{g*gygbgugvgZfzgXftgqgrgogTdmgngcgYfpgfgLfagVf4eybEbCbXd7dSf,f>fNf;etcTfWfRfUfPf>fJfQfHfOfFfKfMfIf?fifDfGfBfEf\\\\}f-fCf@fAf|f*f.f?dhfffGe2e1atc1aobwcubwble,b9dIdge6e9efeff\\\\{frezffe1bldwb+byeZdVb8b1bEbxb;a:bfe6a@d1d5ePa:eqemcZaWeQehc5b-are0d-ctbldyewbwe3bxb,b;a<bfe:breaeye8bEc,bxb2b2btb;a?aWd7e>dmereoe7dpdfeEbYdHafe-e-eFaGakexb-bFc4a-afe.b\\\\{b+cMajaPanePcfe@dIdeeGa+bxd9dSdPabeGa5a@dSd3bDbBb9d>dHd@dobIdRaYaOaVafbVaib9dob>d6d4d-a?a;a>a-aPaBaxc7dVaNaUa?a?a1d1d-aebcb/a1dxcvbpbEaVc7bBaEaBaFa@anb+btbub.b+bzb>bMaHbNc5a1b3b2bDc2b>b:bpb?aDaCa;a;a=anb-!![2iba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"o3j[2|pa\\\\})3(f\\\\{#(tnirP;)R3F*cbVc|b-aWbybHa/axc-bxcGb:aIaDblc:avb|b+bub4bcb-b.c,c*cHaQbJaGaxbNb-b8a1bxbwbtbxbUa-b.b|b3bvbxbfbucsc3bHaHbtcsb/atcobJaub:b6a5aDbtb,b-awb|b.bibHa7bxbzbxbeb-a3b1b.b/b,b|bHaebdb-a,btb1bzb.b1bAbob5a3b-b|b1b/b/a5aJa2bt6Aka721(f\\\\{#,43i7Bja8361(f\\\\{# D4[O31da512Q3a::[R34ma1714(f\\\\{#q\\\\})4;6c:6[O32da88996[R38ea9946j:[O;?ba&[2iha=s,y=z,Y4[\\\\}:2da327-8[O=9da519-8[-8?haq\\\\})6984:6[%89da9418?[YD[D4[YDtca42t8[XD:ca939?o=6[vC2ba5EFH>6Nca72l:[1?Bea420496[R3:ca63d<F1?[D4[D4,ca45[BGt8Oba42FalLkyay,]99999[gnirtS wen=][c n3aea\\\\{)v]y3b&a(niam diov citats cilbup\\\\{RQ ssalc17[w9[D4[/7oca38v9[E4:ca08GW[(ICca0696[(I:ca30j:[HWG8a cdln&&&&;maertStnirP/oi/avajL tuo/metsyS/g"));
$write("%s",("nal/avaj2>b&ategn&&&&2 kcats timil.n&&&&]; V);o?a;3ecaL[\\\\{?av?hha dohtem;3a/4nga repus~3acaRQ83cgassalc.X6[-:2ca79#D[-::ca14!$Ka-:[D43ca30DP[w8;ca538A[E5Bca07wVa96[O?6ba6%T[8ACoa(=:s;0=:c=:i;),@ajaerudecorph5[O32ca69+Ea88[D[5da14588[ZYBda236-N[N?;ca77C?[AS[D4[hErca51gP[s8:ca32:=ara&(tnirp.biL.oken\\\\{D?bianoitcnuf\\\\{Mb/Y[H8[D4[O3wda823H8[<A9ca90bIaRJ[O4>ca5996[95:ca45j:[m>8ca10D4a06[?A5mPbqa(rtStup=niam\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'tni.L[5?=kawohsn\\\\})291cIFi<Mca1488[:5:ba2<5a.6[;52da228i<[;5:da454/6[a[8ba99?[?=<ga4(f\\\\{#=DF[-A>~?b&a(amirpmi oicDAx\\\\})6904(f\\\\{#3Cx\\\\})631d7[R3:wa692(f\\\\{#ni;RQ omtiroglag7[\\\\}G2I6bL5aea.tmf(Rcfacnuf;Y4[Y49datmfE4[E4:raropmi;niam egakca|I[lB4ca02?8dbap/8[I4:ba-C4[C49jatnirp \"\"),\"& VbLf &\"(\"\"tesK4[xI3ba0:Paban/P[VC7*a15(f\\\\{#(,s(llAetirW"));
$write("%s",(";)(resUtxeTtuptuO=:P6[p>3ba5@8fG4[G48daS CE4[O39ca&(C4[.68ba x8[x8[E4[O3\\\\{iaRQ margo76[O3;jaS D : ; R>6[O3:ba\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'C4[O39qa. EPYT B C : ; AR4[;6:ka)*,*(ETIRWM4[E6;haA B : ;K4[O39ba [2cJ4[;6<ba:G4Is[Cga(f\\\\{#(>\\\\{MBba3hOabafiOFba5aPa\\\\{aetirwf:oin\\\\})8(f\\\\{#>-)_(niamp3cL6Bka(f\\\\{# cnirpPIBb6a,atnirP\\\\{)(niaM diov\\\\{noitacilppA:RQ ssalc[\\\\{7B%6ew4aram diov;oidts.dts d[ar4?kaenil-etirw~6|ca(,%3\\\\{cas%G3|nagol.elosnoc;)n5?[2.h4lxa nioj.)1+n(yarrA>-)n(=fd6\\\\{ia!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}54,1\\\\{.v3kja# qes-er(.5lba&?5.ba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"u6\\\\{D3|#3.h40la1% ecalper.-6|z7l[Cntarts(# pam(]YALPSID\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&3kta.NOISIVID ERUDECORP&4\\\\{ma.RQ .DI-MARG23#j4doaNOITACIFITNEDI+3kra[tac-yzal(s[qesodX5c\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'a!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}\\\\}!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");return 0;\\\\}/****/e3a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");s=\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";while 0<len(d):\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\n x as int,y as int=d;i=3;if(n=(x-5)%92+(y-5)%92*87)>3999:\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\n  for _ in range(((d[2]cast int-5)%92+6)):s+=s[len(s)+4000-n]\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\n else:s+=d[2:i=n+2]\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\n d=d[i:]\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\na=0;for i in range(len(s)):b as int=s[i];a-=b;print((\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'*-a if 0>a else\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'-\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'*a)+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\');a=b\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");gsub(/!/,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",s);for(print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"define void f(n)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";for(m=128;m;m/=2)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\""));
$write("%s",("\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,4,:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";if(n/m%2<1)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\};\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"389**6+44*6+00p29*,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";++j<=length(s);print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"f(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"n\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")for(n=9;substr(s,j,1)!=sprintf(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"%c\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",++n););print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,@\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nquit\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")');\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"J\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+a)OD\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\"\");end;\\\"\")\\nsys.exit 0}\"\")]]></xsl:template>"));
$write("%s",("</xsl:stylesheet>\":s=\"   \":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:Console.Write(s &n &Chr(9)&n &\"  \"):Next:Console.Write(n &n &n):End Sub:End Module"));
end endmodule